

module victim_cache(
    input logic clk,
    input logic rst

    
);




logic [255:0] data [8];





endmodule : victim_cache

 